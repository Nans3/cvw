calseab@rivendell.ecen.okstate.edu.7336:1706287626