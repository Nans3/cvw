calseab@rivendell.ecen.okstate.edu.7141:1706287626